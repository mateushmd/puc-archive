/*
	Guia_0304.v
	842536 - Mateus Henrique Medeiros Diniz
*/

module Guia_0304;
	reg [15 : 0] n1 [0 : 4];
	reg [15 : 0] n2 [0 : 4];
	reg [15 : 0] ans;
	
	initial
	begin: main
		n1[0] = 'b11001;
		n1[1] = 'b101_1101;
		n1[2] = 'b110110;
		n1[3] = 'o376;
		n1[4] = 'h7d2;
		
		n2[0] = 'b1101;
		n2[1] = 'b10_0100;
		n2[2] = 'b101101;
		n2[3] = 'o267;
		n2[4] = 'ha51;
				
		$write("a) %b - %b = ", n1[0], n2[0]);
		
		n2[0] = ~n2[0];
		n2[0] = n2[0] + 1;
		ans = n1[0] + n2[0];
		
		$write("%b\n", ans);
		
		$write("b) %b.%b - %b.%b = ", n1[1][6 : 4], n1[1][3 : 0], n2[1][5 : 4], n2[1][3 : 0]);
		
		n2[1] = ~n2[1];
		n2[1] = n2[1] + 1;
		ans = n1[1] + n2[1];
		
		$write("%b.%b\n", ans[6 : 4], ans[3 : 0]);
		
		$write("c) %b - %b = ", n1[2], n2[2]);
		
		n2[2] = ~n2[2];
		n2[2] = n2[2] + 1;
		ans = n1[2] + n2[2];
		
		$write("%b%b\n", ans[3 : 2], ans[1 : 0]);
		
		$write("d) %o - %o = ", n1[3], n2[3]);
		
		n2[3] = ~n2[3];
		n2[3] = n2[3] + 1;
		ans = n1[3] + n2[3];
		
		$write("%o\n", ans);
		
		$write("e) %h - %h = ", n1[4], n2[4]);
		
		n2[4] = ~n2[4];
		n2[4] = n2[4] + 1;
		ans = n1[4] + n2[4];
		
		$write("-%h\n", ans[11 : 0]);
	end
endmodule

/*
	Saída:
	
	a) 0000000000011001 - 0000000000001101 = 0000000000001100
	b) 101.1101 - 10.0100 = 011.1001
	c) 0000000000110110 - 0000000000101101 = 1001
	d) 000376 - 000267 = 000107
	e) 07d2 - 0a51 = -d81
*/